// Verilog
// c2670
// Ninputs 233
// Noutputs 140
// NtotalGates 1269
// BUFF1 272
// AND2 203
// NOT1 321
// AND4 11
// AND3 112
// NAND2 254
// OR2 51
// OR4 22
// NOR2 12
// AND5 7
// OR3 2
// OR5 2

module c2670 (N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
              N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
              N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
              N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
              N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
              N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
              N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
              N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
              N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
              N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
              N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
              N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
              N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
              N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
              N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
              N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
              N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
              N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
              N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
              N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
              N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
              N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
              N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
              N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,
              N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,
              N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,
              N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
              N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,
              N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,
              N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,
              N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,
              N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,
              N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,
              N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,
              N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,
              N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
              N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,
              N216_O,N217_O,N218_O);

input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
      N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
      N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
      N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
      N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
      N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
      N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
      N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
      N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
      N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
      N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
      N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
      N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
      N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
      N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
      N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
      N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
      N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
      N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
      N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
      N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
      N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
      N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
      N216_I,N217_I,N218_I;

output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,
       N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
       N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,
       N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
       N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,
       N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
       N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,
       N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
       N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,
       N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
       N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,
       N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
       N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,
       N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;

wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,
     N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,
     N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,
     N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,
     N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,
     N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,
     N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,
     N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
     N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,
     N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,
     N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,
     N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,
     N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,
     N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,
     N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
     N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,
     N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,
     N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,
     N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
     N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
     N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
     N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
     N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
     N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
     N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
     N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,
     N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
     N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,
     N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,
     N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
     N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,
     N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,
     N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,
     N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,
     N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
     N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
     N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,
     N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
     N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,
     N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,
     N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,
     N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,
     N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,
     N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,
     N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,
     N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
     N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
     N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
     N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
     N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,
     N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,
     N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,
     N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,
     N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
     N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,
     N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,
     N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,
     N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,
     N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,
     N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,
     N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,
     N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
     N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
     N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,
     N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,
     N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,
     N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,
     N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,
     N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,
     N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
     N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,
     N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
     N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,
     N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,
     N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,
     N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,
     N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,
     N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
     N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
     N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,
     N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,
     N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,
     N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,
     N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,
     N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,
     N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
     N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,
     N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,
     N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,
     N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,
     N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,
     N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,
     N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
     N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
     N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
     N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,
     N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,
     N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,
     N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,
     N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,
     N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,
     N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
     N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,
     N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,
     N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,
     N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,
     N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,
     N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
     N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
     N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877,N4000,N4001,N4002;

buf BUFF1_1 (N398, N219);
buf BUFF1_2 (N400, N219);
buf BUFF1_3 (N401, N219);
and AND2_4 (N405, N1, N3);
not NOT1_5 (N408, N230);
buf BUFF1_6 (N419, N253);
buf BUFF1_7 (N420, N253);
not NOT1_8 (N425, N262);
buf BUFF1_9 (N456, N290);
buf BUFF1_10 (N457, N290);
buf BUFF1_11 (N458, N290);
and AND4_12 (N485, N309, N305, N301, N297);
not NOT1_13 (N486, N405);
not NOT1_14 (N487, N44);
not NOT1_15 (N488, N132);
not NOT1_16 (N489, N82);
not NOT1_17 (N490, N96);
not NOT1_18 (N491, N69);
not NOT1_19 (N492, N120);
not NOT1_20 (N493, N57);
not NOT1_21 (N494, N108);
and AND3_22 (N495, N2, N15, N237);
buf BUFF1_23 (N496, N237);
and AND2_24 (N499, N37, N37);
buf BUFF1_25 (N500, N219);
buf BUFF1_26 (N503, N8);
buf BUFF1_27 (N506, N8);
buf BUFF1_28 (N509, N227);
buf BUFF1_29 (N521, N234);
not NOT1_30 (N533, N241);
not NOT1_31 (N537, N246);
and AND2_32 (N543, N11, N246);
and AND4_33 (N544, N132, N82, N96, N44);
and AND4_34 (N547, N120, N57, N108, N69);
buf BUFF1_35 (N550, N227);
buf BUFF1_36 (N562, N234);
not NOT1_37 (N574, N256);
not NOT1_38 (N578, N259);
buf BUFF1_39 (N582, N319);
buf BUFF1_40 (N594, N322);
not NOT1_41 (N606, N328);
not NOT1_42 (N607, N331);
not NOT1_43 (N608, N334);
not NOT1_44 (N609, N337);
not NOT1_45 (N610, N340);
not NOT1_46 (N611, N343);
not NOT1_47 (N612, N352);
buf BUFF1_48 (N613, N319);
buf BUFF1_49 (N625, N322);
buf BUFF1_50 (N637, N16);
buf BUFF1_51 (N643, N16);
not NOT1_52 (N650, N355);
and AND2_53 (N651, N7, N237);
not NOT1_54 (N655, N263);
not NOT1_55 (N659, N266);
not NOT1_56 (N663, N269);
not NOT1_57 (N667, N272);
not NOT1_58 (N671, N275);
not NOT1_59 (N675, N278);
not NOT1_60 (N679, N281);
not NOT1_61 (N683, N284);
not NOT1_62 (N687, N287);
buf BUFF1_63 (N693, N29);
buf BUFF1_64 (N699, N29);
not NOT1_65 (N705, N294);
not NOT1_66 (N711, N297);
not NOT1_67 (N715, N301);
not NOT1_68 (N719, N305);
not NOT1_69 (N723, N309);
not NOT1_70 (N727, N313);
not NOT1_71 (N730, N316);
not NOT1_72 (N733, N346);
not NOT1_73 (N734, N349);
buf BUFF1_74 (N735, N259);
buf BUFF1_75 (N738, N256);
buf BUFF1_76 (N741, N263);
buf BUFF1_77 (N744, N269);
buf BUFF1_78 (N747, N266);
buf BUFF1_79 (N750, N275);
buf BUFF1_80 (N753, N272);
buf BUFF1_81 (N756, N281);
buf BUFF1_82 (N759, N278);
buf BUFF1_83 (N762, N287);
buf BUFF1_84 (N765, N284);
buf BUFF1_85 (N768, N294);
buf BUFF1_86 (N771, N301);
buf BUFF1_87 (N774, N297);
buf BUFF1_88 (N777, N309);
buf BUFF1_89 (N780, N305);
buf BUFF1_90 (N783, N316);
buf BUFF1_91 (N786, N313);
not NOT1_92 (N792, N485);
not NOT1_93 (N799, N495);
not NOT1_94 (N800, N499);
buf BUFF1_95 (N805, N500);
nand NAND2_96 (N900, N331, N606);
nand NAND2_97 (N901, N328, N607);
nand NAND2_98 (N902, N337, N608);
nand NAND2_99 (N903, N334, N609);
nand NAND2_100 (N904, N343, N610);
nand NAND2_101 (N905, N340, N611);
nand NAND2_102 (N998, N349, N733);
nand NAND2_103 (N999, N346, N734);
and AND2_104 (N1026, N94, N500);
and AND2_105 (N1027, N325, N651);
not NOT1_106 (N1028, N651);
nand NAND2_107 (N1029, N231, N651);
not NOT1_108 (N1032, N544);
not NOT1_109 (N1033, N547);
and AND2_110 (N1034, N547, N544);
buf BUFF1_111 (N1037, N503);
not NOT1_112 (N1042, N509);
not NOT1_113 (N1053, N521);
and AND3_114 (N1064, N80, N509, N521);
and AND3_115 (N1065, N68, N509, N521);
and AND3_116 (N1066, N79, N509, N521);
and AND3_117 (N1067, N78, N509, N521);
and AND3_118 (N1068, N77, N509, N521);
and AND2_119 (N1069, N11, N537);
buf BUFF1_120 (N1070, N503);
not NOT1_121 (N1075, N550);
not NOT1_122 (N1086, N562);
and AND3_123 (N1097, N76, N550, N562);
and AND3_124 (N1098, N75, N550, N562);
and AND3_125 (N1099, N74, N550, N562);
and AND3_126 (N1100, N73, N550, N562);
and AND3_127 (N1101, N72, N550, N562);
not NOT1_128 (N1102, N582);
not NOT1_129 (N1113, N594);
and AND3_130 (N1124, N114, N582, N594);
and AND3_131 (N1125, N113, N582, N594);
and AND3_132 (N1126, N112, N582, N594);
and AND3_133 (N1127, N111, N582, N594);
and AND2_134 (N1128, N582, N594);
nand NAND2_135 (N1129, N900, N901);
nand NAND2_136 (N1133, N902, N903);
nand NAND2_137 (N1137, N904, N905);
not NOT1_138 (N1140, N741);
nand NAND2_139 (N1141, N741, N612);
not NOT1_140 (N1142, N744);
not NOT1_141 (N1143, N747);
not NOT1_142 (N1144, N750);
not NOT1_143 (N1145, N753);
not NOT1_144 (N1146, N613);
not NOT1_145 (N1157, N625);
and AND3_146 (N1168, N118, N613, N625);
and AND3_147 (N1169, N107, N613, N625);
and AND3_148 (N1170, N117, N613, N625);
and AND3_149 (N1171, N116, N613, N625);
and AND3_150 (N1172, N115, N613, N625);
not NOT1_151 (N1173, N637);
not NOT1_152 (N1178, N643);
not NOT1_153 (N1184, N768);
nand NAND2_154 (N1185, N768, N650);
not NOT1_155 (N1186, N771);
not NOT1_156 (N1187, N774);
not NOT1_157 (N1188, N777);
not NOT1_158 (N1189, N780);
buf BUFF1_159 (N1190, N506);
buf BUFF1_160 (N1195, N506);
not NOT1_161 (N1200, N693);
not NOT1_162 (N1205, N699);
not NOT1_163 (N1210, N735);
not NOT1_164 (N1211, N738);
not NOT1_165 (N1212, N756);
not NOT1_166 (N1213, N759);
not NOT1_167 (N1214, N762);
not NOT1_168 (N1215, N765);
nand NAND2_169 (N1216, N998, N999);
buf BUFF1_170 (N1219, N574);
buf BUFF1_171 (N1222, N578);
buf BUFF1_172 (N1225, N655);
buf BUFF1_173 (N1228, N659);
buf BUFF1_174 (N1231, N663);
buf BUFF1_175 (N1234, N667);
buf BUFF1_176 (N1237, N671);
buf BUFF1_177 (N1240, N675);
buf BUFF1_178 (N1243, N679);
buf BUFF1_179 (N1246, N683);
not NOT1_180 (N1249, N783);
not NOT1_181 (N1250, N786);
buf BUFF1_182 (N1251, N687);
buf BUFF1_183 (N1254, N705);
buf BUFF1_184 (N1257, N711);
buf BUFF1_185 (N1260, N715);
buf BUFF1_186 (N1263, N719);
buf BUFF1_187 (N1266, N723);
not NOT1_188 (N1269, N1027);
and AND2_189 (N1275, N325, N1032);
and AND2_190 (N1276, N231, N1033);
buf BUFF1_191 (N1277, N1034);
or OR2_192 (N1302, N1069, N543);
nand NAND2_193 (N1351, N352, N1140);
nand NAND2_194 (N1352, N747, N1142);
nand NAND2_195 (N1353, N744, N1143);
nand NAND2_196 (N1354, N753, N1144);
nand NAND2_197 (N1355, N750, N1145);
nand NAND2_198 (N1395, N355, N1184);
nand NAND2_199 (N1396, N774, N1186);
nand NAND2_200 (N1397, N771, N1187);
nand NAND2_201 (N1398, N780, N1188);
nand NAND2_202 (N1399, N777, N1189);
nand NAND2_203 (N1422, N738, N1210);
nand NAND2_204 (N1423, N735, N1211);
nand NAND2_205 (N1424, N759, N1212);
nand NAND2_206 (N1425, N756, N1213);
nand NAND2_207 (N1426, N765, N1214);
nand NAND2_208 (N1427, N762, N1215);
nand NAND2_209 (N1440, N786, N1249);
nand NAND2_210 (N1441, N783, N1250);
not NOT1_211 (N1448, N1034);
not NOT1_212 (N1449, N1275);
not NOT1_213 (N1450, N1276);
and AND3_214 (N1451, N93, N1042, N1053);
and AND3_215 (N1452, N55, N509, N1053);
and AND3_216 (N1453, N67, N1042, N521);
and AND3_217 (N1454, N81, N1042, N1053);
and AND3_218 (N1455, N43, N509, N1053);
and AND3_219 (N1456, N56, N1042, N521);
and AND3_220 (N1457, N92, N1042, N1053);
and AND3_221 (N1458, N54, N509, N1053);
and AND3_222 (N1459, N66, N1042, N521);
and AND3_223 (N1460, N91, N1042, N1053);
and AND3_224 (N1461, N53, N509, N1053);
and AND3_225 (N1462, N65, N1042, N521);
and AND3_226 (N1463, N90, N1042, N1053);
and AND3_227 (N1464, N52, N509, N1053);
and AND3_228 (N1465, N64, N1042, N521);
and AND3_229 (N1466, N89, N1075, N1086);
and AND3_230 (N1467, N51, N550, N1086);
and AND3_231 (N1468, N63, N1075, N562);
and AND3_232 (N1469, N88, N1075, N1086);
and AND3_233 (N1470, N50, N550, N1086);
and AND3_234 (N1471, N62, N1075, N562);
and AND3_235 (N1472, N87, N1075, N1086);
and AND3_236 (N1473, N49, N550, N1086);
and AND2_237 (N1474, N1075, N562);
and AND3_238 (N1475, N86, N1075, N1086);
and AND3_239 (N1476, N48, N550, N1086);
and AND3_240 (N1477, N61, N1075, N562);
and AND3_241 (N1478, N85, N1075, N1086);
and AND3_242 (N1479, N47, N550, N1086);
and AND3_243 (N1480, N60, N1075, N562);
and AND3_244 (N1481, N138, N1102, N1113);
and AND3_245 (N1482, N102, N582, N1113);
and AND3_246 (N1483, N126, N1102, N594);
and AND3_247 (N1484, N137, N1102, N1113);
and AND3_248 (N1485, N101, N582, N1113);
and AND3_249 (N1486, N125, N1102, N594);
and AND3_250 (N1487, N136, N1102, N1113);
and AND3_251 (N1488, N100, N582, N1113);
and AND3_252 (N1489, N124, N1102, N594);
and AND3_253 (N1490, N135, N1102, N1113);
and AND3_254 (N1491, N99, N582, N1113);
and AND3_255 (N1492, N123, N1102, N594);
and AND2_256 (N1493, N1102, N1113);
and AND2_257 (N1494, N582, N1113);
and AND2_258 (N1495, N1102, N594);
not NOT1_259 (N1496, N1129);
not NOT1_260 (N1499, N1133);
nand NAND2_261 (N1502, N1351, N1141);
nand NAND2_262 (N1506, N1352, N1353);
nand NAND2_263 (N1510, N1354, N1355);
buf BUFF1_264 (N1513, N1137);
buf BUFF1_265 (N1516, N1137);
not NOT1_266 (N1519, N1219);
not NOT1_267 (N1520, N1222);
not NOT1_268 (N1521, N1225);
not NOT1_269 (N1522, N1228);
not NOT1_270 (N1523, N1231);
not NOT1_271 (N1524, N1234);
not NOT1_272 (N1525, N1237);
not NOT1_273 (N1526, N1240);
not NOT1_274 (N1527, N1243);
not NOT1_275 (N1528, N1246);
and AND3_276 (N1529, N142, N1146, N1157);
and AND3_277 (N1530, N106, N613, N1157);
and AND3_278 (N1531, N130, N1146, N625);
and AND3_279 (N1532, N131, N1146, N1157);
and AND3_280 (N1533, N95, N613, N1157);
and AND3_281 (N1534, N119, N1146, N625);
and AND3_282 (N1535, N141, N1146, N1157);
and AND3_283 (N1536, N105, N613, N1157);
and AND3_284 (N1537, N129, N1146, N625);
and AND3_285 (N1538, N140, N1146, N1157);
and AND3_286 (N1539, N104, N613, N1157);
and AND3_287 (N1540, N128, N1146, N625);
and AND3_288 (N1541, N139, N1146, N1157);
and AND3_289 (N1542, N103, N613, N1157);
and AND3_290 (N1543, N127, N1146, N625);
and AND2_291 (N1544, N19, N1173);
and AND2_292 (N1545, N4, N1173);
and AND2_293 (N1546, N20, N1173);
and AND2_294 (N1547, N5, N1173);
and AND2_295 (N1548, N21, N1178);
and AND2_296 (N1549, N22, N1178);
and AND2_297 (N1550, N23, N1178);
and AND2_298 (N1551, N6, N1178);
and AND2_299 (N1552, N24, N1178);
nand NAND2_300 (N1553, N1395, N1185);
nand NAND2_301 (N1557, N1396, N1397);
nand NAND2_302 (N1561, N1398, N1399);
and AND2_303 (N1564, N25, N1200);
and AND2_304 (N1565, N32, N1200);
and AND2_305 (N1566, N26, N1200);
and AND2_306 (N1567, N33, N1200);
and AND2_307 (N1568, N27, N1205);
and AND2_308 (N1569, N34, N1205);
and AND2_309 (N1570, N35, N1205);
and AND2_310 (N1571, N28, N1205);
not NOT1_311 (N1572, N1251);
not NOT1_312 (N1573, N1254);
not NOT1_313 (N1574, N1257);
not NOT1_314 (N1575, N1260);
not NOT1_315 (N1576, N1263);
not NOT1_316 (N1577, N1266);
nand NAND2_317 (N1578, N1422, N1423);
not NOT1_318 (N1581, N1216);
nand NAND2_319 (N1582, N1426, N1427);
nand NAND2_320 (N1585, N1424, N1425);
nand NAND2_321 (N1588, N1440, N1441);
and AND2_322 (N1591, N1449, N1450);
or OR4_323 (N1596, N1451, N1452, N1453, N1064);
or OR4_324 (N1600, N1454, N1455, N1456, N1065);
or OR4_325 (N1606, N1457, N1458, N1459, N1066);
or OR4_326 (N1612, N1460, N1461, N1462, N1067);
or OR4_327 (N1615, N1463, N1464, N1465, N1068);
or OR4_328 (N1619, N1466, N1467, N1468, N1097);
or OR4_329 (N1624, N1469, N1470, N1471, N1098);
or OR4_330 (N1628, N1472, N1473, N1474, N1099);
or OR4_331 (N1631, N1475, N1476, N1477, N1100);
or OR4_332 (N1634, N1478, N1479, N1480, N1101);
or OR4_333 (N1637, N1481, N1482, N1483, N1124);
or OR4_334 (N1642, N1484, N1485, N1486, N1125);
or OR4_335 (N1647, N1487, N1488, N1489, N1126);
or OR4_336 (N1651, N1490, N1491, N1492, N1127);
or OR4_337 (N1656, N1493, N1494, N1495, N1128);
or OR4_338 (N1676, N1532, N1533, N1534, N1169);
or OR4_339 (N1681, N1535, N1536, N1537, N1170);
or OR4_340 (N1686, N1538, N1539, N1540, N1171);
or OR4_341 (N1690, N1541, N1542, N1543, N1172);
or OR4_342 (N1708, N1529, N1530, N1531, N1168);
buf BUFF1_343 (N1726, N1591);
not NOT1_344 (N1770, N1502);
not NOT1_345 (N1773, N1506);
not NOT1_346 (N1776, N1513);
not NOT1_347 (N1777, N1516);
buf BUFF1_348 (N1778, N1510);
buf BUFF1_349 (N1781, N1510);
and AND3_350 (N1784, N1133, N1129, N1513);
and AND3_351 (N1785, N1499, N1496, N1516);
not NOT1_352 (N1795, N1553);
not NOT1_353 (N1798, N1557);
buf BUFF1_354 (N1801, N1561);
buf BUFF1_355 (N1804, N1561);
not NOT1_356 (N1807, N1588);
not NOT1_357 (N1808, N1578);
nand NAND2_358 (N1809, N1578, N1581);
not NOT1_359 (N1810, N1582);
not NOT1_360 (N1811, N1585);
and AND2_361 (N1813, N1596, N241);
and AND2_362 (N1814, N1606, N241);
and AND2_363 (N1815, N1600, N241);
not NOT1_364 (N1816, N1642);
not NOT1_365 (N1817, N1647);
not NOT1_366 (N1818, N1637);
not NOT1_367 (N1819, N1624);
not NOT1_368 (N1820, N1619);
not NOT1_369 (N1821, N1615);
and AND4_370 (N1822, N496, N224, N36, N1591);
and AND4_371 (N1823, N496, N224, N1591, N486);
buf BUFF1_372 (N1824, N1596);
not NOT1_373 (N1827, N1606);
and AND2_374 (N1830, N1600, N537);
and AND2_375 (N1831, N1606, N537);
and AND2_376 (N1832, N1619, N246);
not NOT1_377 (N1833, N1596);
not NOT1_378 (N1836, N1600);
not NOT1_379 (N1841, N1606);
buf BUFF1_380 (N1848, N1612);
buf BUFF1_381 (N1852, N1615);
buf BUFF1_382 (N1856, N1619);
buf BUFF1_383 (N1863, N1624);
buf BUFF1_384 (N1870, N1628);
buf BUFF1_385 (N1875, N1631);
buf BUFF1_386 (N1880, N1634);
nand NAND2_387 (N1885, N727, N1651);
nand NAND2_388 (N1888, N730, N1656);
buf BUFF1_389 (N1891, N1686);
and AND2_390 (N1894, N1637, N425);
not NOT1_391 (N1897, N1642);
and AND3_392 (N1908, N1496, N1133, N1776);
and AND3_393 (N1909, N1129, N1499, N1777);
and AND2_394 (N1910, N1600, N637);
and AND2_395 (N1911, N1606, N637);
and AND2_396 (N1912, N1612, N637);
and AND2_397 (N1913, N1615, N637);
and AND2_398 (N1914, N1619, N643);
and AND2_399 (N1915, N1624, N643);
and AND2_400 (N1916, N1628, N643);
and AND2_401 (N1917, N1631, N643);
and AND2_402 (N1918, N1634, N643);
not NOT1_403 (N1919, N1708);
and AND2_404 (N1928, N1676, N693);
and AND2_405 (N1929, N1681, N693);
and AND2_406 (N1930, N1686, N693);
and AND2_407 (N1931, N1690, N693);
and AND2_408 (N1932, N1637, N699);
and AND2_409 (N1933, N1642, N699);
and AND2_410 (N1934, N1647, N699);
and AND2_411 (N1935, N1651, N699);
buf BUFF1_412 (N1936, N1600);
nand NAND2_413 (N1939, N1216, N1808);
nand NAND2_414 (N1940, N1585, N1810);
nand NAND2_415 (N1941, N1582, N1811);
buf BUFF1_416 (N1942, N1676);
buf BUFF1_417 (N1945, N1686);
buf BUFF1_418 (N1948, N1681);
buf BUFF1_419 (N1951, N1637);
buf BUFF1_420 (N1954, N1690);
buf BUFF1_421 (N1957, N1647);
buf BUFF1_422 (N1960, N1642);
buf BUFF1_423 (N1963, N1656);
buf BUFF1_424 (N1966, N1651);
or OR2_425 (N1969, N533, N1815);
not NOT1_426 (N1970, N1822);
not NOT1_427 (N1971, N1823);
buf BUFF1_428 (N2010, N1848);
buf BUFF1_429 (N2012, N1852);
buf BUFF1_430 (N2014, N1856);
buf BUFF1_431 (N2016, N1863);
buf BUFF1_432 (N2018, N1870);
buf BUFF1_433 (N2020, N1875);
buf BUFF1_434 (N2022, N1880);
not NOT1_435 (N2028, N1778);
not NOT1_436 (N2029, N1781);
nor NOR2_437 (N2030, N1908, N1784);
nor NOR2_438 (N2031, N1909, N1785);
and AND3_439 (N2032, N1506, N1502, N1778);
and AND3_440 (N2033, N1773, N1770, N1781);
or OR2_441 (N2034, N1571, N1935);
not NOT1_442 (N2040, N1801);
not NOT1_443 (N2041, N1804);
and AND3_444 (N2042, N1557, N1553, N1801);
and AND3_445 (N2043, N1798, N1795, N1804);
nand NAND2_446 (N2046, N1939, N1809);
nand NAND2_447 (N2049, N1940, N1941);
or OR2_448 (N2052, N1544, N1910);
or OR2_449 (N2055, N1545, N1911);
or OR2_450 (N2058, N1546, N1912);
or OR2_451 (N2061, N1547, N1913);
or OR2_452 (N2064, N1548, N1914);
or OR2_453 (N2067, N1549, N1915);
or OR2_454 (N2070, N1550, N1916);
or OR2_455 (N2073, N1551, N1917);
or OR2_456 (N2076, N1552, N1918);
or OR2_457 (N2079, N1564, N1928);
or OR2_458 (N2095, N1565, N1929);
or OR2_459 (N2098, N1566, N1930);
or OR2_460 (N2101, N1567, N1931);
or OR2_461 (N2104, N1568, N1932);
or OR2_462 (N2107, N1569, N1933);
or OR2_463 (N2110, N1570, N1934);
and AND3_464 (N2113, N1897, N1894, N40);
not NOT1_465 (N2119, N1894);
nand NAND2_466 (N2120, N408, N1827);
and AND2_467 (N2125, N1824, N537);
and AND2_468 (N2126, N1852, N246);
and AND2_469 (N2127, N1848, N537);
not NOT1_470 (N2128, N1848);
not NOT1_471 (N2135, N1852);
not NOT1_472 (N2141, N1863);
not NOT1_473 (N2144, N1870);
not NOT1_474 (N2147, N1875);
not NOT1_475 (N2150, N1880);
and AND2_476 (N2153, N727, N1885);
and AND2_477 (N2154, N1885, N1651);
and AND2_478 (N2155, N730, N1888);
and AND2_479 (N2156, N1888, N1656);
and AND3_480 (N2157, N1770, N1506, N2028);
and AND3_481 (N2158, N1502, N1773, N2029);
not NOT1_482 (N2171, N1942);
nand NAND2_483 (N2172, N1942, N1919);
not NOT1_484 (N2173, N1945);
not NOT1_485 (N2174, N1948);
not NOT1_486 (N2175, N1951);
not NOT1_487 (N2176, N1954);
and AND3_488 (N2177, N1795, N1557, N2040);
and AND3_489 (N2178, N1553, N1798, N2041);
buf BUFF1_490 (N2185, N1836);
buf BUFF1_491 (N2188, N1833);
buf BUFF1_492 (N2191, N1841);
not NOT1_493 (N2194, N1856);
not NOT1_494 (N2197, N1827);
not NOT1_495 (N2200, N1936);
buf BUFF1_496 (N2201, N1836);
buf BUFF1_497 (N2204, N1833);
buf BUFF1_498 (N2207, N1841);
buf BUFF1_499 (N2210, N1824);
buf BUFF1_500 (N2213, N1841);
buf BUFF1_501 (N2216, N1841);
nand NAND2_502 (N2219, N2031, N2030);
not NOT1_503 (N2234, N1957);
not NOT1_504 (N2235, N1960);
not NOT1_505 (N2236, N1963);
not NOT1_506 (N2237, N1966);
and AND3_507 (N2250, N40, N1897, N2119);
or OR2_508 (N2266, N1831, N2126);
or OR2_509 (N2269, N2127, N1832);
or OR2_510 (N2291, N2153, N2154);
or OR2_511 (N2294, N2155, N2156);
nor NOR2_512 (N2297, N2157, N2032);
nor NOR2_513 (N2298, N2158, N2033);
not NOT1_514 (N2300, N2046);
not NOT1_515 (N2301, N2049);
nand NAND2_516 (N2302, N2052, N1519);
not NOT1_517 (N2303, N2052);
nand NAND2_518 (N2304, N2055, N1520);
not NOT1_519 (N2305, N2055);
nand NAND2_520 (N2306, N2058, N1521);
not NOT1_521 (N2307, N2058);
nand NAND2_522 (N2308, N2061, N1522);
not NOT1_523 (N2309, N2061);
nand NAND2_524 (N2310, N2064, N1523);
not NOT1_525 (N2311, N2064);
nand NAND2_526 (N2312, N2067, N1524);
not NOT1_527 (N2313, N2067);
nand NAND2_528 (N2314, N2070, N1525);
not NOT1_529 (N2315, N2070);
nand NAND2_530 (N2316, N2073, N1526);
not NOT1_531 (N2317, N2073);
nand NAND2_532 (N2318, N2076, N1527);
not NOT1_533 (N2319, N2076);
nand NAND2_534 (N2320, N2079, N1528);
not NOT1_535 (N2321, N2079);
nand NAND2_536 (N2322, N1708, N2171);
nand NAND2_537 (N2323, N1948, N2173);
nand NAND2_538 (N2324, N1945, N2174);
nand NAND2_539 (N2325, N1954, N2175);
nand NAND2_540 (N2326, N1951, N2176);
nor NOR2_541 (N2327, N2177, N2042);
nor NOR2_542 (N2328, N2178, N2043);
nand NAND2_543 (N2329, N2095, N1572);
not NOT1_544 (N2330, N2095);
nand NAND2_545 (N2331, N2098, N1573);
not NOT1_546 (N2332, N2098);
nand NAND2_547 (N2333, N2101, N1574);
not NOT1_548 (N2334, N2101);
nand NAND2_549 (N2335, N2104, N1575);
not NOT1_550 (N2336, N2104);
nand NAND2_551 (N2337, N2107, N1576);
not NOT1_552 (N2338, N2107);
nand NAND2_553 (N2339, N2110, N1577);
not NOT1_554 (N2340, N2110);
nand NAND2_555 (N2354, N1960, N2234);
nand NAND2_556 (N2355, N1957, N2235);
nand NAND2_557 (N2356, N1966, N2236);
nand NAND2_558 (N2357, N1963, N2237);
and AND2_559 (N2358, N2120, N533);
not NOT1_560 (N2359, N2113);
not NOT1_561 (N2364, N2185);
not NOT1_562 (N2365, N2188);
not NOT1_563 (N2366, N2191);
not NOT1_564 (N2367, N2194);
buf BUFF1_565 (N2368, N2120);
not NOT1_566 (N2372, N2201);
not NOT1_567 (N2373, N2204);
not NOT1_568 (N2374, N2207);
not NOT1_569 (N2375, N2210);
not NOT1_570 (N2376, N2213);
not NOT1_571 (N2377, N2113);
buf BUFF1_572 (N2382, N2113);
and AND2_573 (N2386, N2120, N246);
buf BUFF1_574 (N2387, N2266);
buf BUFF1_575 (N2388, N2266);
buf BUFF1_576 (N2389, N2269);
buf BUFF1_577 (N2390, N2269);
buf BUFF1_578 (N2391, N2113);
not NOT1_579 (N2395, N2113);
nand NAND2_580 (N2400, N2219, N2300);
not NOT1_581 (N2403, N2216);
not NOT1_582 (N2406, N2219);
nand NAND2_583 (N2407, N1219, N2303);
nand NAND2_584 (N2408, N1222, N2305);
nand NAND2_585 (N2409, N1225, N2307);
nand NAND2_586 (N2410, N1228, N2309);
nand NAND2_587 (N2411, N1231, N2311);
nand NAND2_588 (N2412, N1234, N2313);
nand NAND2_589 (N2413, N1237, N2315);
nand NAND2_590 (N2414, N1240, N2317);
nand NAND2_591 (N2415, N1243, N2319);
nand NAND2_592 (N2416, N1246, N2321);
nand NAND2_593 (N2417, N2322, N2172);
nand NAND2_594 (N2421, N2323, N2324);
nand NAND2_595 (N2425, N2325, N2326);
nand NAND2_596 (N2428, N1251, N2330);
nand NAND2_597 (N2429, N1254, N2332);
nand NAND2_598 (N2430, N1257, N2334);
nand NAND2_599 (N2431, N1260, N2336);
nand NAND2_600 (N2432, N1263, N2338);
nand NAND2_601 (N2433, N1266, N2340);
buf BUFF1_602 (N2434, N2128);
buf BUFF1_603 (N2437, N2135);
buf BUFF1_604 (N2440, N2144);
buf BUFF1_605 (N2443, N2141);
buf BUFF1_606 (N2446, N2150);
buf BUFF1_607 (N2449, N2147);
not NOT1_608 (N2452, N2197);
nand NAND2_609 (N2453, N2197, N2200);
buf BUFF1_610 (N2454, N2128);
buf BUFF1_611 (N2457, N2144);
buf BUFF1_612 (N2460, N2141);
buf BUFF1_613 (N2463, N2150);
buf BUFF1_614 (N2466, N2147);
not NOT1_615 (N2469, N2120);
buf BUFF1_616 (N2472, N2128);
buf BUFF1_617 (N2475, N2135);
buf BUFF1_618 (N2478, N2128);
buf BUFF1_619 (N2481, N2135);
nand NAND2_620 (N2484, N2298, N2297);
nand NAND2_621 (N2487, N2356, N2357);
nand NAND2_622 (N2490, N2354, N2355);
nand NAND2_623 (N2493, N2328, N2327);
or OR2_624 (N2496, N2358, N1814);
nand NAND2_625 (N2503, N2188, N2364);
nand NAND2_626 (N2504, N2185, N2365);
nand NAND2_627 (N2510, N2204, N2372);
nand NAND2_628 (N2511, N2201, N2373);
or OR2_629 (N2521, N1830, N2386);
nand NAND2_630 (N2528, N2046, N2406);
not NOT1_631 (N2531, N2291);
not NOT1_632 (N2534, N2294);
buf BUFF1_633 (N2537, N2250);
buf BUFF1_634 (N2540, N2250);
nand NAND2_635 (N2544, N2302, N2407);
nand NAND2_636 (N2545, N2304, N2408);
nand NAND2_637 (N2546, N2306, N2409);
nand NAND2_638 (N2547, N2308, N2410);
nand NAND2_639 (N2548, N2310, N2411);
nand NAND2_640 (N2549, N2312, N2412);
nand NAND2_641 (N2550, N2314, N2413);
nand NAND2_642 (N2551, N2316, N2414);
nand NAND2_643 (N2552, N2318, N2415);
nand NAND2_644 (N2553, N2320, N2416);
nand NAND2_645 (N2563, N2329, N2428);
nand NAND2_646 (N2564, N2331, N2429);
nand NAND2_647 (N2565, N2333, N2430);
nand NAND2_648 (N2566, N2335, N2431);
nand NAND2_649 (N2567, N2337, N2432);
nand NAND2_650 (N2568, N2339, N2433);
nand NAND2_651 (N2579, N1936, N2452);
buf BUFF1_652 (N2603, N2359);
and AND2_653 (N2607, N1880, N2377);
and AND2_654 (N2608, N1676, N2377);
and AND2_655 (N2609, N1681, N2377);
and AND2_656 (N2610, N1891, N2377);
and AND2_657 (N2611, N1856, N2382);
and AND2_658 (N2612, N1863, N2382);
nand NAND2_659 (N2613, N2503, N2504);
not NOT1_660 (N2617, N2434);
nand NAND2_661 (N2618, N2434, N2366);
nand NAND2_662 (N2619, N2437, N2367);
not NOT1_663 (N2620, N2437);
not NOT1_664 (N2621, N2368);
nand NAND2_665 (N2624, N2510, N2511);
not NOT1_666 (N2628, N2454);
nand NAND2_667 (N2629, N2454, N2374);
not NOT1_668 (N2630, N2472);
and AND2_669 (N2631, N1856, N2391);
and AND2_670 (N2632, N1863, N2391);
and AND2_671 (N2633, N1880, N2395);
and AND2_672 (N2634, N1676, N2395);
and AND2_673 (N2635, N1681, N2395);
and AND2_674 (N2636, N1891, N2395);
not NOT1_675 (N2638, N2382);
buf BUFF1_676 (N2643, N2521);
buf BUFF1_677 (N2644, N2521);
not NOT1_678 (N2645, N2475);
not NOT1_679 (N2646, N2391);
nand NAND2_680 (N2652, N2528, N2400);
not NOT1_681 (N2655, N2478);
not NOT1_682 (N2656, N2481);
buf BUFF1_683 (N2659, N2359);
not NOT1_684 (N2663, N2484);
nand NAND2_685 (N2664, N2484, N2301);
not NOT1_686 (N2665, N2553);
not NOT1_687 (N2666, N2552);
not NOT1_688 (N2667, N2551);
not NOT1_689 (N2668, N2550);
not NOT1_690 (N2669, N2549);
not NOT1_691 (N2670, N2548);
not NOT1_692 (N2671, N2547);
not NOT1_693 (N2672, N2546);
not NOT1_694 (N2673, N2545);
not NOT1_695 (N2674, N2544);
not NOT1_696 (N2675, N2568);
not NOT1_697 (N2676, N2567);
not NOT1_698 (N2677, N2566);
not NOT1_699 (N2678, N2565);
not NOT1_700 (N2679, N2564);
not NOT1_701 (N2680, N2563);
not NOT1_702 (N2681, N2417);
not NOT1_703 (N2684, N2421);
buf BUFF1_704 (N2687, N2425);
buf BUFF1_705 (N2690, N2425);
not NOT1_706 (N2693, N2493);
nand NAND2_707 (N2694, N2493, N1807);
not NOT1_708 (N2695, N2440);
not NOT1_709 (N2696, N2443);
not NOT1_710 (N2697, N2446);
not NOT1_711 (N2698, N2449);
not NOT1_712 (N2699, N2457);
not NOT1_713 (N2700, N2460);
not NOT1_714 (N2701, N2463);
not NOT1_715 (N2702, N2466);
nand NAND2_716 (N2703, N2579, N2453);
not NOT1_717 (N2706, N2469);
not NOT1_718 (N2707, N2487);
not NOT1_719 (N2708, N2490);
and AND2_720 (N2709, N2294, N2534);
and AND2_721 (N2710, N2291, N2531);
nand NAND2_722 (N2719, N2191, N2617);
nand NAND2_723 (N2720, N2194, N2620);
nand NAND2_724 (N2726, N2207, N2628);
buf BUFF1_725 (N2729, N2537);
buf BUFF1_726 (N2738, N2537);
not NOT1_727 (N2743, N2652);
nand NAND2_728 (N2747, N2049, N2663);
and AND5_729 (N2748, N2665, N2666, N2667, N2668, N2669);
and AND5_730 (N2749, N2670, N2671, N2672, N2673, N2674);
and AND2_731 (N2750, N2034, N2675);
and AND5_732 (N2751, N2676, N2677, N2678, N2679, N2680);
nand NAND2_733 (N2760, N1588, N2693);
buf BUFF1_734 (N2761, N2540);
buf BUFF1_735 (N2766, N2540);
nand NAND2_736 (N2771, N2443, N2695);
nand NAND2_737 (N2772, N2440, N2696);
nand NAND2_738 (N2773, N2449, N2697);
nand NAND2_739 (N2774, N2446, N2698);
nand NAND2_740 (N2775, N2460, N2699);
nand NAND2_741 (N2776, N2457, N2700);
nand NAND2_742 (N2777, N2466, N2701);
nand NAND2_743 (N2778, N2463, N2702);
nand NAND2_744 (N2781, N2490, N2707);
nand NAND2_745 (N2782, N2487, N2708);
or OR2_746 (N2783, N2709, N2534);
or OR2_747 (N2784, N2710, N2531);
and AND2_748 (N2789, N1856, N2638);
and AND2_749 (N2790, N1863, N2638);
and AND2_750 (N2791, N1870, N2638);
and AND2_751 (N2792, N1875, N2638);
not NOT1_752 (N2793, N2613);
nand NAND2_753 (N2796, N2719, N2618);
nand NAND2_754 (N2800, N2619, N2720);
not NOT1_755 (N2803, N2624);
nand NAND2_756 (N2806, N2726, N2629);
and AND2_757 (N2809, N1856, N2646);
and AND2_758 (N2810, N1863, N2646);
and AND2_759 (N2811, N1870, N2646);
and AND2_760 (N2812, N1875, N2646);
and AND2_761 (N2817, N2743, N14);
buf BUFF1_762 (N2820, N2603);
nand NAND2_763 (N2826, N2747, N2664);
and AND2_764 (N2829, N2748, N2749);
and AND2_765 (N2830, N2750, N2751);
buf BUFF1_766 (N2831, N2659);
not NOT1_767 (N2837, N2687);
not NOT1_768 (N2838, N2690);
and AND3_769 (N2839, N2421, N2417, N2687);
and AND3_770 (N2840, N2684, N2681, N2690);
nand NAND2_771 (N2841, N2760, N2694);
buf BUFF1_772 (N2844, N2603);
buf BUFF1_773 (N2854, N2603);
buf BUFF1_774 (N2859, N2659);
buf BUFF1_775 (N2869, N2659);
nand NAND2_776 (N2874, N2773, N2774);
nand NAND2_777 (N2877, N2771, N2772);
not NOT1_778 (N2880, N2703);
nand NAND2_779 (N2881, N2703, N2706);
nand NAND2_780 (N2882, N2777, N2778);
nand NAND2_781 (N2885, N2775, N2776);
nand NAND2_782 (N2888, N2781, N2782);
nand NAND2_783 (N2891, N2783, N2784);
and AND2_784 (N2894, N2607, N2729);
and AND2_785 (N2895, N2608, N2729);
and AND2_786 (N2896, N2609, N2729);
and AND2_787 (N2897, N2610, N2729);
or OR2_788 (N2898, N2789, N2611);
or OR2_789 (N2899, N2790, N2612);
and AND2_790 (N2900, N2791, N1037);
and AND2_791 (N2901, N2792, N1037);
or OR2_792 (N2914, N2809, N2631);
or OR2_793 (N2915, N2810, N2632);
and AND2_794 (N2916, N2811, N1070);
and AND2_795 (N2917, N2812, N1070);
and AND2_796 (N2918, N2633, N2738);
and AND2_797 (N2919, N2634, N2738);
and AND2_798 (N2920, N2635, N2738);
and AND2_799 (N2921, N2636, N2738);
buf BUFF1_800 (N2925, N2817);
and AND3_801 (N2931, N2829, N2830, N1302);
and AND3_802 (N2938, N2681, N2421, N2837);
and AND3_803 (N2939, N2417, N2684, N2838);
nand NAND2_804 (N2963, N2469, N2880);
not NOT1_805 (N2970, N2841);
not NOT1_806 (N2971, N2826);
not NOT1_807 (N2972, N2894);
not NOT1_808 (N2975, N2895);
not NOT1_809 (N2978, N2896);
not NOT1_810 (N2981, N2897);
and AND2_811 (N2984, N2898, N1037);
and AND2_812 (N2985, N2899, N1037);
not NOT1_813 (N2986, N2900);
not NOT1_814 (N2989, N2901);
not NOT1_815 (N2992, N2796);
buf BUFF1_816 (N2995, N2800);
buf BUFF1_817 (N2998, N2800);
buf BUFF1_818 (N3001, N2806);
buf BUFF1_819 (N3004, N2806);
and AND2_820 (N3007, N574, N2820);
and AND2_821 (N3008, N2914, N1070);
and AND2_822 (N3009, N2915, N1070);
not NOT1_823 (N3010, N2916);
not NOT1_824 (N3013, N2917);
not NOT1_825 (N3016, N2918);
not NOT1_826 (N3019, N2919);
not NOT1_827 (N3022, N2920);
not NOT1_828 (N3025, N2921);
not NOT1_829 (N3028, N2817);
and AND2_830 (N3029, N574, N2831);
not NOT1_831 (N3030, N2820);
and AND2_832 (N3035, N578, N2820);
and AND2_833 (N3036, N655, N2820);
and AND2_834 (N3037, N659, N2820);
buf BUFF1_835 (N3038, N2931);
not NOT1_836 (N3039, N2831);
and AND2_837 (N3044, N578, N2831);
and AND2_838 (N3045, N655, N2831);
and AND2_839 (N3046, N659, N2831);
nor NOR2_840 (N3047, N2938, N2839);
nor NOR2_841 (N3048, N2939, N2840);
not NOT1_842 (N3049, N2888);
not NOT1_843 (N3050, N2844);
and AND2_844 (N3053, N663, N2844);
and AND2_845 (N3054, N667, N2844);
and AND2_846 (N3055, N671, N2844);
and AND2_847 (N3056, N675, N2844);
and AND2_848 (N3057, N679, N2854);
and AND2_849 (N3058, N683, N2854);
and AND2_850 (N3059, N687, N2854);
and AND2_851 (N3060, N705, N2854);
not NOT1_852 (N3061, N2859);
and AND2_853 (N3064, N663, N2859);
and AND2_854 (N3065, N667, N2859);
and AND2_855 (N3066, N671, N2859);
and AND2_856 (N3067, N675, N2859);
and AND2_857 (N3068, N679, N2869);
and AND2_858 (N3069, N683, N2869);
and AND2_859 (N3070, N687, N2869);
and AND2_860 (N3071, N705, N2869);
not NOT1_861 (N3072, N2874);
not NOT1_862 (N3073, N2877);
not NOT1_863 (N3074, N2882);
not NOT1_864 (N3075, N2885);
nand NAND2_865 (N3076, N2881, N2963);
not NOT1_866 (N3079, N2931);
not NOT1_867 (N3088, N2984);
not NOT1_868 (N3091, N2985);
not NOT1_869 (N3110, N3008);
not NOT1_870 (N3113, N3009);
and AND2_871 (N3137, N3055, N1190);
and AND2_872 (N3140, N3056, N1190);
and AND2_873 (N3143, N3057, N2761);
and AND2_874 (N3146, N3058, N2761);
and AND2_875 (N3149, N3059, N2761);
and AND2_876 (N3152, N3060, N2761);
and AND2_877 (N3157, N3066, N1195);
and AND2_878 (N3160, N3067, N1195);
and AND2_879 (N3163, N3068, N2766);
and AND2_880 (N3166, N3069, N2766);
and AND2_881 (N3169, N3070, N2766);
and AND2_882 (N3172, N3071, N2766);
nand NAND2_883 (N3175, N2877, N3072);
nand NAND2_884 (N3176, N2874, N3073);
nand NAND2_885 (N3177, N2885, N3074);
nand NAND2_886 (N3178, N2882, N3075);
nand NAND2_887 (N3180, N3048, N3047);
not NOT1_888 (N3187, N2995);
not NOT1_889 (N3188, N2998);
not NOT1_890 (N3189, N3001);
not NOT1_891 (N3190, N3004);
and AND3_892 (N3191, N2796, N2613, N2995);
and AND3_893 (N3192, N2992, N2793, N2998);
and AND3_894 (N3193, N2624, N2368, N3001);
and AND3_895 (N3194, N2803, N2621, N3004);
nand NAND2_896 (N3195, N3076, N2375);
not NOT1_897 (N3196, N3076);
and AND2_898 (N3197, N687, N3030);
and AND2_899 (N3208, N687, N3039);
and AND2_900 (N3215, N705, N3030);
and AND2_901 (N3216, N711, N3030);
and AND2_902 (N3217, N715, N3030);
and AND2_903 (N3218, N705, N3039);
and AND2_904 (N3219, N711, N3039);
and AND2_905 (N3220, N715, N3039);
and AND2_906 (N3222, N719, N3050);
and AND2_907 (N3223, N723, N3050);
and AND2_908 (N3230, N719, N3061);
and AND2_909 (N3231, N723, N3061);
nand NAND2_910 (N3238, N3175, N3176);
nand NAND2_911 (N3241, N3177, N3178);
buf BUFF1_912 (N3244, N2981);
buf BUFF1_913 (N3247, N2978);
buf BUFF1_914 (N3250, N2975);
buf BUFF1_915 (N3253, N2972);
buf BUFF1_916 (N3256, N2989);
buf BUFF1_917 (N3259, N2986);
buf BUFF1_918 (N3262, N3025);
buf BUFF1_919 (N3265, N3022);
buf BUFF1_920 (N3268, N3019);
buf BUFF1_921 (N3271, N3016);
buf BUFF1_922 (N3274, N3013);
buf BUFF1_923 (N3277, N3010);
and AND3_924 (N3281, N2793, N2796, N3187);
and AND3_925 (N3282, N2613, N2992, N3188);
and AND3_926 (N3283, N2621, N2624, N3189);
and AND3_927 (N3284, N2368, N2803, N3190);
nand NAND2_928 (N3286, N2210, N3196);
or OR2_929 (N3288, N3197, N3007);
nand NAND2_930 (N3289, N3180, N3049);
and AND2_931 (N3291, N3152, N2981);
and AND2_932 (N3293, N3149, N2978);
and AND2_933 (N3295, N3146, N2975);
and AND2_934 (N3296, N2972, N3143);
and AND2_935 (N3299, N3140, N2989);
and AND2_936 (N3301, N3137, N2986);
or OR2_937 (N3302, N3208, N3029);
and AND2_938 (N3304, N3172, N3025);
and AND2_939 (N3306, N3169, N3022);
and AND2_940 (N3308, N3166, N3019);
and AND2_941 (N3309, N3016, N3163);
and AND2_942 (N3312, N3160, N3013);
and AND2_943 (N3314, N3157, N3010);
or OR2_944 (N3315, N3215, N3035);
or OR2_945 (N3318, N3216, N3036);
or OR2_946 (N3321, N3217, N3037);
or OR2_947 (N3324, N3218, N3044);
or OR2_948 (N3327, N3219, N3045);
or OR2_949 (N3330, N3220, N3046);
not NOT1_950 (N3333, N3180);
or OR2_951 (N3334, N3222, N3053);
or OR2_952 (N3335, N3223, N3054);
or OR2_953 (N3336, N3230, N3064);
or OR2_954 (N3337, N3231, N3065);
buf BUFF1_955 (N3340, N3152);
buf BUFF1_956 (N3344, N3149);
buf BUFF1_957 (N3348, N3146);
buf BUFF1_958 (N3352, N3143);
buf BUFF1_959 (N3356, N3140);
buf BUFF1_960 (N3360, N3137);
buf BUFF1_961 (N3364, N3091);
buf BUFF1_962 (N3367, N3088);
buf BUFF1_963 (N3370, N3172);
buf BUFF1_964 (N3374, N3169);
buf BUFF1_965 (N3378, N3166);
buf BUFF1_966 (N3382, N3163);
buf BUFF1_967 (N3386, N3160);
buf BUFF1_968 (N3390, N3157);
buf BUFF1_969 (N3394, N3113);
buf BUFF1_970 (N3397, N3110);
nand NAND2_971 (N3400, N3195, N3286);
nor NOR2_972 (N3401, N3281, N3191);
nor NOR2_973 (N3402, N3282, N3192);
nor NOR2_974 (N3403, N3283, N3193);
nor NOR2_975 (N3404, N3284, N3194);
not NOT1_976 (N3405, N3238);
not NOT1_977 (N3406, N3241);
and AND2_978 (N3409, N3288, N1836);
nand NAND2_979 (N3410, N2888, N3333);
not NOT1_980 (N3412, N3244);
not NOT1_981 (N3414, N3247);
not NOT1_982 (N3416, N3250);
not NOT1_983 (N3418, N3253);
not NOT1_984 (N3420, N3256);
not NOT1_985 (N3422, N3259);
and AND2_986 (N3428, N3302, N1836);
not NOT1_987 (N3430, N3262);
not NOT1_988 (N3432, N3265);
not NOT1_989 (N3434, N3268);
not NOT1_990 (N3436, N3271);
not NOT1_991 (N3438, N3274);
not NOT1_992 (N3440, N3277);
and AND2_993 (N3450, N3334, N1190);
and AND2_994 (N3453, N3335, N1190);
and AND2_995 (N3456, N3336, N1195);
and AND2_996 (N3459, N3337, N1195);
and AND2_997 (N3478, N3400, N533);
and AND2_998 (N3479, N3318, N2128);
and AND2_999 (N3480, N3315, N1841);
nand NAND2_1000 (N3481, N3410, N3289);
not NOT1_1001 (N3482, N3340);
nand NAND2_1002 (N3483, N3340, N3412);
not NOT1_1003 (N3484, N3344);
nand NAND2_1004 (N3485, N3344, N3414);
not NOT1_1005 (N3486, N3348);
nand NAND2_1006 (N3487, N3348, N3416);
not NOT1_1007 (N3488, N3352);
nand NAND2_1008 (N3489, N3352, N3418);
not NOT1_1009 (N3490, N3356);
nand NAND2_1010 (N3491, N3356, N3420);
not NOT1_1011 (N3492, N3360);
nand NAND2_1012 (N3493, N3360, N3422);
not NOT1_1013 (N3494, N3364);
not NOT1_1014 (N3496, N3367);
and AND2_1015 (N3498, N3321, N2135);
and AND2_1016 (N3499, N3327, N2128);
and AND2_1017 (N3500, N3324, N1841);
not NOT1_1018 (N3501, N3370);
nand NAND2_1019 (N3502, N3370, N3430);
not NOT1_1020 (N3503, N3374);
nand NAND2_1021 (N3504, N3374, N3432);
not NOT1_1022 (N3505, N3378);
nand NAND2_1023 (N3506, N3378, N3434);
not NOT1_1024 (N3507, N3382);
nand NAND2_1025 (N3508, N3382, N3436);
not NOT1_1026 (N3509, N3386);
nand NAND2_1027 (N3510, N3386, N3438);
not NOT1_1028 (N3511, N3390);
nand NAND2_1029 (N3512, N3390, N3440);
not NOT1_1030 (N3513, N3394);
not NOT1_1031 (N3515, N3397);
and AND2_1032 (N3517, N3330, N2135);
nand NAND2_1033 (N3522, N3402, N3401);
nand NAND2_1034 (N3525, N3404, N3403);
buf BUFF1_1035 (N3528, N3318);
buf BUFF1_1036 (N3531, N3315);
buf BUFF1_1037 (N3534, N3321);
buf BUFF1_1038 (N3537, N3327);
buf BUFF1_1039 (N3540, N3324);
buf BUFF1_1040 (N3543, N3330);
or OR2_1041 (N3546, N3478, N1813);
not NOT1_1042 (N3551, N3481);
nand NAND2_1043 (N3552, N3244, N3482);
nand NAND2_1044 (N3553, N3247, N3484);
nand NAND2_1045 (N3554, N3250, N3486);
nand NAND2_1046 (N3555, N3253, N3488);
nand NAND2_1047 (N3556, N3256, N3490);
nand NAND2_1048 (N3557, N3259, N3492);
and AND2_1049 (N3558, N3453, N3091);
and AND2_1050 (N3559, N3450, N3088);
nand NAND2_1051 (N3563, N3262, N3501);
nand NAND2_1052 (N3564, N3265, N3503);
nand NAND2_1053 (N3565, N3268, N3505);
nand NAND2_1054 (N3566, N3271, N3507);
nand NAND2_1055 (N3567, N3274, N3509);
nand NAND2_1056 (N3568, N3277, N3511);
and AND2_1057 (N3569, N3459, N3113);
and AND2_1058 (N3570, N3456, N3110);
buf BUFF1_1059 (N3576, N3453);
buf BUFF1_1060 (N3579, N3450);
buf BUFF1_1061 (N3585, N3459);
buf BUFF1_1062 (N3588, N3456);
not NOT1_1063 (N3592, N3522);
nand NAND2_1064 (N3593, N3522, N3405);
not NOT1_1065 (N3594, N3525);
nand NAND2_1066 (N3595, N3525, N3406);
not NOT1_1067 (N3596, N3528);
nand NAND2_1068 (N3597, N3528, N2630);
nand NAND2_1069 (N3598, N3531, N2376);
not NOT1_1070 (N3599, N3531);
and AND2_1071 (N3600, N3551, N800);
nand NAND2_1072 (N3603, N3552, N3483);
nand NAND2_1073 (N3608, N3553, N3485);
nand NAND2_1074 (N3612, N3554, N3487);
nand NAND2_1075 (N3615, N3555, N3489);
nand NAND2_1076 (N3616, N3556, N3491);
nand NAND2_1077 (N3622, N3557, N3493);
not NOT1_1078 (N3629, N3534);
nand NAND2_1079 (N3630, N3534, N2645);
not NOT1_1080 (N3631, N3537);
nand NAND2_1081 (N3632, N3537, N2655);
nand NAND2_1082 (N3633, N3540, N2403);
not NOT1_1083 (N3634, N3540);
nand NAND2_1084 (N3635, N3563, N3502);
nand NAND2_1085 (N3640, N3564, N3504);
nand NAND2_1086 (N3644, N3565, N3506);
nand NAND2_1087 (N3647, N3566, N3508);
nand NAND2_1088 (N3648, N3567, N3510);
nand NAND2_1089 (N3654, N3568, N3512);
not NOT1_1090 (N3661, N3543);
nand NAND2_1091 (N3662, N3543, N2656);
nand NAND2_1092 (N3667, N3238, N3592);
nand NAND2_1093 (N3668, N3241, N3594);
nand NAND2_1094 (N3669, N2472, N3596);
nand NAND2_1095 (N3670, N2213, N3599);
buf BUFF1_1096 (N3671, N3600);
not NOT1_1097 (N3691, N3576);
nand NAND2_1098 (N3692, N3576, N3494);
not NOT1_1099 (N3693, N3579);
nand NAND2_1100 (N3694, N3579, N3496);
nand NAND2_1101 (N3695, N2475, N3629);
nand NAND2_1102 (N3696, N2478, N3631);
nand NAND2_1103 (N3697, N2216, N3634);
not NOT1_1104 (N3716, N3585);
nand NAND2_1105 (N3717, N3585, N3513);
not NOT1_1106 (N3718, N3588);
nand NAND2_1107 (N3719, N3588, N3515);
nand NAND2_1108 (N3720, N2481, N3661);
nand NAND2_1109 (N3721, N3667, N3593);
nand NAND2_1110 (N3722, N3668, N3595);
nand NAND2_1111 (N3723, N3669, N3597);
nand NAND2_1112 (N3726, N3670, N3598);
not NOT1_1113 (N3727, N3600);
nand NAND2_1114 (N3728, N3364, N3691);
nand NAND2_1115 (N3729, N3367, N3693);
nand NAND2_1116 (N3730, N3695, N3630);
and AND4_1117 (N3731, N3608, N3615, N3612, N3603);
not NOT1_1 (N4000, N3731);
xor XOR2_1 (N4001, N3731, N4000);
or OR2_1 (N4002, N4000, N4001);
and AND2_1118 (N3732, N3603, N3293);
and AND3_1119 (N3733, N3608, N3603, N3295);
and AND4_1120 (N3734, N3612, N3603, N3296, N3608);
and AND2_1121 (N3735, N3616, N3301);
and AND3_1122 (N3736, N3622, N3616, N3558);
nand NAND2_1123 (N3737, N3696, N3632);
nand NAND2_1124 (N3740, N3697, N3633);
nand NAND2_1125 (N3741, N3394, N3716);
nand NAND2_1126 (N3742, N3397, N3718);
nand NAND2_1127 (N3743, N3720, N3662);
and AND4_1128 (N3744, N3640, N3647, N3644, N3635);
and AND2_1129 (N3745, N3635, N3306);
and AND3_1130 (N3746, N3640, N3635, N3308);
and AND4_1131 (N3747, N3644, N3635, N3309, N3640);
and AND2_1132 (N3748, N3648, N3314);
and AND3_1133 (N3749, N3654, N3648, N3569);
not NOT1_1134 (N3750, N3721);
and AND2_1135 (N3753, N3722, N246);
nand NAND2_1136 (N3754, N3728, N3692);
nand NAND2_1137 (N3758, N3729, N3694);
not NOT1_1138 (N3761, N4002);
or OR4_1139 (N3762, N3291, N3732, N3733, N3734);
nand NAND2_1140 (N3767, N3741, N3717);
nand NAND2_1141 (N3771, N3742, N3719);
not NOT1_1142 (N3774, N3744);
or OR4_1143 (N3775, N3304, N3745, N3746, N3747);
and AND2_1144 (N3778, N3723, N3480);
and AND3_1145 (N3779, N3726, N3723, N3409);
or OR2_1146 (N3780, N2125, N3753);
and AND2_1147 (N3790, N3750, N800);
and AND2_1148 (N3793, N3737, N3500);
and AND3_1149 (N3794, N3740, N3737, N3428);
or OR3_1150 (N3802, N3479, N3778, N3779);
buf BUFF1_1151 (N3803, N3780);
buf BUFF1_1152 (N3804, N3780);
not NOT1_1153 (N3805, N3762);
and AND5_1154 (N3806, N3622, N3730, N3754, N3616, N3758);
and AND4_1155 (N3807, N3754, N3616, N3559, N3622);
and AND5_1156 (N3808, N3758, N3754, N3616, N3498, N3622);
buf BUFF1_1157 (N3809, N3790);
or OR3_1158 (N3811, N3499, N3793, N3794);
not NOT1_1159 (N3812, N3775);
and AND5_1160 (N3813, N3654, N3743, N3767, N3648, N3771);
and AND4_1161 (N3814, N3767, N3648, N3570, N3654);
and AND5_1162 (N3815, N3771, N3767, N3648, N3517, N3654);
or OR5_1163 (N3816, N3299, N3735, N3736, N3807, N3808);
and AND2_1164 (N3817, N3806, N3802);
nand NAND2_1165 (N3818, N3805, N3761);
not NOT1_1166 (N3819, N3790);
or OR5_1167 (N3820, N3312, N3748, N3749, N3814, N3815);
and AND2_1168 (N3821, N3813, N3811);
nand NAND2_1169 (N3822, N3812, N3774);
or OR2_1170 (N3823, N3816, N3817);
and AND3_1171 (N3826, N3727, N3819, N2841);
or OR2_1172 (N3827, N3820, N3821);
not NOT1_1173 (N3834, N3823);
and AND2_1174 (N3835, N3818, N3823);
not NOT1_1175 (N3836, N3827);
and AND2_1176 (N3837, N3822, N3827);
and AND2_1177 (N3838, N3762, N3834);
and AND2_1178 (N3839, N3775, N3836);
or OR2_1179 (N3840, N3838, N3835);
or OR2_1180 (N3843, N3839, N3837);
buf BUFF1_1181 (N3851, N3843);
nand NAND2_1182 (N3852, N3843, N3840);
and AND2_1183 (N3857, N3843, N3852);
and AND2_1184 (N3858, N3852, N3840);
or OR2_1185 (N3859, N3857, N3858);
not NOT1_1186 (N3864, N3859);
and AND2_1187 (N3869, N3859, N3864);
or OR2_1188 (N3870, N3869, N3864);
not NOT1_1189 (N3875, N3870);
and AND3_1190 (N3876, N2826, N3028, N3870);
and AND3_1191 (N3877, N3826, N3876, N1591);
buf BUFF1_1192 (N3881, N3877);
not NOT1_1193 (N3882, N3877);
buf BUFF1_1194 (N143_O, N143_I);
buf BUFF1_1195 (N144_O, N144_I);
buf BUFF1_1196 (N145_O, N145_I);
buf BUFF1_1197 (N146_O, N146_I);
buf BUFF1_1198 (N147_O, N147_I);
buf BUFF1_1199 (N148_O, N148_I);
buf BUFF1_1200 (N149_O, N149_I);
buf BUFF1_1201 (N150_O, N150_I);
buf BUFF1_1202 (N151_O, N151_I);
buf BUFF1_1203 (N152_O, N152_I);
buf BUFF1_1204 (N153_O, N153_I);
buf BUFF1_1205 (N154_O, N154_I);
buf BUFF1_1206 (N155_O, N155_I);
buf BUFF1_1207 (N156_O, N156_I);
buf BUFF1_1208 (N157_O, N157_I);
buf BUFF1_1209 (N158_O, N158_I);
buf BUFF1_1210 (N159_O, N159_I);
buf BUFF1_1211 (N160_O, N160_I);
buf BUFF1_1212 (N161_O, N161_I);
buf BUFF1_1213 (N162_O, N162_I);
buf BUFF1_1214 (N163_O, N163_I);
buf BUFF1_1215 (N164_O, N164_I);
buf BUFF1_1216 (N165_O, N165_I);
buf BUFF1_1217 (N166_O, N166_I);
buf BUFF1_1218 (N167_O, N167_I);
buf BUFF1_1219 (N168_O, N168_I);
buf BUFF1_1220 (N169_O, N169_I);
buf BUFF1_1221 (N170_O, N170_I);
buf BUFF1_1222 (N171_O, N171_I);
buf BUFF1_1223 (N172_O, N172_I);
buf BUFF1_1224 (N173_O, N173_I);
buf BUFF1_1225 (N174_O, N174_I);
buf BUFF1_1226 (N175_O, N175_I);
buf BUFF1_1227 (N176_O, N176_I);
buf BUFF1_1228 (N177_O, N177_I);
buf BUFF1_1229 (N178_O, N178_I);
buf BUFF1_1230 (N179_O, N179_I);
buf BUFF1_1231 (N180_O, N180_I);
buf BUFF1_1232 (N181_O, N181_I);
buf BUFF1_1233 (N182_O, N182_I);
buf BUFF1_1234 (N183_O, N183_I);
buf BUFF1_1235 (N184_O, N184_I);
buf BUFF1_1236 (N185_O, N185_I);
buf BUFF1_1237 (N186_O, N186_I);
buf BUFF1_1238 (N187_O, N187_I);
buf BUFF1_1239 (N188_O, N188_I);
buf BUFF1_1240 (N189_O, N189_I);
buf BUFF1_1241 (N190_O, N190_I);
buf BUFF1_1242 (N191_O, N191_I);
buf BUFF1_1243 (N192_O, N192_I);
buf BUFF1_1244 (N193_O, N193_I);
buf BUFF1_1245 (N194_O, N194_I);
buf BUFF1_1246 (N195_O, N195_I);
buf BUFF1_1247 (N196_O, N196_I);
buf BUFF1_1248 (N197_O, N197_I);
buf BUFF1_1249 (N198_O, N198_I);
buf BUFF1_1250 (N199_O, N199_I);
buf BUFF1_1251 (N200_O, N200_I);
buf BUFF1_1252 (N201_O, N201_I);
buf BUFF1_1253 (N202_O, N202_I);
buf BUFF1_1254 (N203_O, N203_I);
buf BUFF1_1255 (N204_O, N204_I);
buf BUFF1_1256 (N205_O, N205_I);
buf BUFF1_1257 (N206_O, N206_I);
buf BUFF1_1258 (N207_O, N207_I);
buf BUFF1_1259 (N208_O, N208_I);
buf BUFF1_1260 (N209_O, N209_I);
buf BUFF1_1261 (N210_O, N210_I);
buf BUFF1_1262 (N211_O, N211_I);
buf BUFF1_1263 (N212_O, N212_I);
buf BUFF1_1264 (N213_O, N213_I);
buf BUFF1_1265 (N214_O, N214_I);
buf BUFF1_1266 (N215_O, N215_I);
buf BUFF1_1267 (N216_O, N216_I);
buf BUFF1_1268 (N217_O, N217_I);
buf BUFF1_1269 (N218_O, N218_I);

endmodule